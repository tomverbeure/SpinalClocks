// Generator : SpinalHDL v1.1.5    git head : 0310b2489a097f2b9de5535e02192d9ddd2764ae
// Date      : 16/12/2018, 23:17:58
// Component : Top


module Top (
      output  io_led_green,
      input   io_switch);
  assign io_led_green = 1'b1;
endmodule

